TestBench2 for Homework3 

Vin 1 0 3
R1 1 2 2k
R1 1 2 a
R1 1 2 2k 123
R1 2 0 100
R2R 2 0 100
C1 2 0 2e-10
L1 2 4 8
.DC Vin 0.5 2 0.1
.Print DC V(2)
.Print wf V(2)
.Print dc V(w)
.Print DC wf V(2)
.end
asf
wfwfwf