TestBench1 for Homework4
* 2022 EDA course testbench netlist
* 2022-10-17

Vin 1 0 3
R1 1 2 200
C1 1 2 20p
R2 2 0 100
L1 2 0 10m

.DC Vin 1 2 0.1
.end    
